`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/17/2024 07:53:02 PM
// Design Name: 
// Module Name: ladder_sprite
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ladder_sprite(
    input logic [5:0] addr,
    output logic [13:0] data
    );
    parameter ADDR_WIDTH = 6;
    parameter DATA_WIDTH = 14;
    parameter [0:49][DATA_WIDTH-1:0] ROM = {
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11111111111111,
    14'b11111111111111,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11111111111111,
    14'b11111111111111,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11111111111111,
    14'b11111111111111,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11111111111111,
    14'b11111111111111,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11111111111111,
    14'b11111111111111,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11111111111111,
    14'b11111111111111,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011,
    14'b11111111111111,
    14'b11111111111111,
    14'b11000000000011,
    14'b11000000000011,
    14'b11000000000011

    };
    
    assign data = ROM[addr];
endmodule
