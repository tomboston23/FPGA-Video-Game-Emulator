`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/18/2024 02:19:55 PM
// Design Name: 
// Module Name: mario_sprite
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mario_sprite(
    input [3:0] X,
    input [3:0] Y,
    output [1:0] pal

    );
    //00 means alpha = 0
    //01 means red
    //10 means dark brown
    //11 means light brown
    
    parameter[0:15][0:31] ROM = {
        32'b00_00_00_00_00_00_00_01_01_01_01_01_01_01_00_00_00_00_00_00,
        32'b00_00_00_00_00_01_01_01_01_01_01_01_01_01_01_01_00_00_00_00,
        32'b00_00_00_10_10_10_10_10_11_11_10_11_00_00_00_00_00_00_00_00,
        32'b00_00_10_10_11_10_11_11_11_11_10_11_11_11_11_10_00_00_00_00,
        32'b00_00_10_10_11_10_10_11_11_11_11_10_11_11_11_11_11_11_00_00,
        32'b00_00_10_10_10_10_11_11_11_11_11_10_10_10_10_10_00_00_00_00,
        32'b00_00_00_00_00_00_11_11_11_11_11_11_11_11_00_00_00_00_00_00,
        32'b00_00_00_00_10_10_10_10_01_10_10_10_10_00_00_00_00_00_00_00,
        32'b00_00_10_10_10_10_01_10_10_10_01_10_10_10_10_00_00_00_00_00,
        32'b00_10_10_10_10_10_01_01_01_01_01_10_10_10_10_10_00_00_00_00,
        32'b00_11_11_11_11_11_10_01_11_10_10_11_01_11_11_00_00_00_00_00,
        32'b00_11_11_11_11_11_10_10_10_10_10_11_11_11_11_11_00_00_00_00,
        32'b00_11_11_11_11_10_10_10_10_10_10_10_11_11_11_11_00_00_00_00,
        32'b00_00_00_00_00_00_01_01_01_01_00_01_01_01_01_01_00_00_00_00,
        32'b00_00_10_10_10_10_00_00_00_00_10_10_10_10_10_00_00_00_00_00,
        32'b00_10_10_10_10_10_00_00_00_00_10_10_10_10_10_10_00_00_00_00
    };
    logic [31:0] data = ROM[Y];
    assign pal = data[X*2 +:2];
    
endmodule
